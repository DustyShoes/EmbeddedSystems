//module child (in, out);
//	input in [3:0];
//	output out [3:0];
//	
//	wire in [3:0];
//	wire out [3:0];
//	
//	//do things
//endmodule
