//module parent (data, returned);
//	input data [3:0];
//	output returned [3:0];
//	wire data [3:0];
//	wire returned [3:0];
//	
//	child ch (
//		.in(data),
//		.out(returned)
//	);
//
//	//do things
//endmodule
