module fulladder3bits(inA, inB, cin, cout, sum);

endmodule
